//////////////////////////////////////////////////////////////////////////////////
//
// top.v
//
// This is the top module of 1-locater within a byte-stream. Consists of two FIFOs
// that at send-in phase respectively store the non-zero inputs and their time to come. 
// At send-out phase, the FIFO is read (while another send-in phase might be running at 
// the same time) and a time span is devoted to each entry depending on its hamming weight. 
// e.g. for 11001011 five clock cycles will be devoted. A decoder, weight_locator, instantly 
// generates the index of ones in that byte. Finally the output location is generated by 
// calculating the time that byte came in (from FIFO2) and the location in byte that the 
// decoder indicates.The input bit-stream is given input_binary.bin which can be 
//
// wrritten by: Morteza Hosseini
//
//////////////////////////////////////////////////////////////////////////////////

`timescale 1ns / 1ps

module top (clk, srst, start, din, hw, locations, valid, overflow);

// Inputs
input clk;//clock
input srst;//reset
input start; // start to send in
input [7:0] din; //data in, which is streamed in the form of an episode of 128 bytes

// Outputs
output reg [7:0] hw; // Hamming Weight. We assign more than 5 bits, to loosen up the computation of hamming weigh in case that FIFO is not yet full
output [9:0] locations; // consecutive locations of 1s from the input at the output. This signal is sent out instantly after din has come in.
output valid; // indicates whether the location is valid. This is essentially used to distinguish a real existing 1 at location=0 from non-existing ones that have a location=0 indicator  
output overflow; // FIFO is limited and is constrained to hold between 31 to 248 1s from each episode (31: one 1 per byte, 248: eight 1s per 31 byte.) Overflow, indicates that FIFO is full

// Wires and Registers
wire rd_en_valid; // this is to lessen the read span with one clock cycle
reg   [7:0] din_reg; // input signals are registered so that a better estimation of reg2reg critical path is given by the CAD tool
reg   start_reg; // input signals are registered so that a better estimation of reg2reg critical path is given by CAD tool
wire  [7:0] hw_read_in; //unlike previous hw, this signal dynamically changes based on any input
reg   [7:0] hw_reg; // We need an accumulator on hamming weights that instantly generates the accumulations with no delay. later at send-out this register is passed to hw output
reg   [7:0] valid_interval; // this reg at the send-out phase counts down as much as the hamming weight in order to indicate the valid span of the output
reg   [7:0] clk_cycle_counter; // this register counts up to indicate at which cycle the state in an episode is 
wire  rd_en; // signal to FIFOs to allow when to read from
wire  wr_en; // signal to FIFOs to allow when to write at
wire  [2:0] location_in_byte; // This signal combines all the 8 signals coming out of the weight_locator an,d by means of 8 mutually exclusive pulses, represent the location of 1s one at a clock cycle
reg   L0_h,L1_h,L2_h,L3_h,L4_h,L5_h,L6_h,L7_h; // These are mutually exclusive pulses that are in fact place holders for the outputs of the weight_locator.

//L0_h__| |___________________
//L1_h____| |_________________
//L2_h______| |_______________
//L3_h________| |_____________
//L4_h__________| |___________
//L5_h____________| |_________
//L6_h_______________| |______
//L7_h_________________| |____

wire  [2:0] L0,L1,L2,L3,L4,L5,L6,L7; // outputs from the weight_locator
reg   rd_en_pulse; // this signal is the first read pulse upon the 128th clock cycle. after this pulse the hamming weigh is passed to the controller and from there on it knows how many more clock cycles to read from the FIFO
wire  [7:0] stored_non_zero_byte; // (stored at first FIFO) non-zero bytes that were saved in FIFO in the read-in phase
wire  [7:0] stored_clk_cycle; // (stored at snd FIFO) time at which the non-zero byte was saved
reg   [3:0] PC_in;	// Hamming weight, A.K.A Population Count, of one single byte in read_in phase
wire  [3:0] PC_out;	// Hamming weight, A.K.A Population Count, of one single byte after sending out
reg   [3:0] PC_out_temp; // PC_out is the instant byte hamming weight value coming from the weight_locator. This PC_out_temp register is the decremental version of PC_out for controlling reasons. (see the signal diagram below this page)

// a Dynamic byte hamming weigh generator at read-in phase. We need this signal to be accumulated to hw_reg
always @(*)
PC_in = din_reg[0]+din_reg[1]+din_reg[2]+din_reg[3]+din_reg[4]+din_reg[5]+din_reg[6]+din_reg[7];

// din_reg: input signals are registered so that a better estimation of reg2reg critical path is given by the CAD tool
always @(posedge clk)
begin
	if (srst==1)
	din_reg <= 0;
	else
	din_reg <= din;
end

// start_reg: input signals are registered so that a better estimation of reg2reg critical path is given by the CAD tool
always @(posedge clk)
begin
	if ((srst==1))
	start_reg <= 0;
	else
	start_reg <= start;
end

// hw_reg: accumulating the weights dynamically in the send-in phase
always @(posedge clk)
begin
	if ((srst==1)||(start_reg==1))
	hw_reg <= 0;
	else if (clk_cycle_counter<128)
	hw_reg <= hw_read_in;
end

// clk_cycle_counter: it resets to zero at the begining of every episode and counts up to 128 (or 255 if un attended by the start signal)
always @(posedge clk)
begin
	if ((srst==1)||(start_reg==1))
	clk_cycle_counter <= 0;
	else
	clk_cycle_counter <= clk_cycle_counter + 1;
end

// valid_interval: a valid interval is equal to the hamming weight of the input. we load it with the hamming weigh, and then it counts down. while it is non-zero we are in valid output region
always @(posedge clk)
begin
  if (clk_cycle_counter == 127)
	valid_interval <= hw_read_in;	
	else if ((srst==1)||(valid_interval<2))
	valid_interval <= 0;
	else 
	valid_interval <= valid_interval - 1;  
end

// hw: hamming weigh, which is sent out, and is latched during the valid interval
always @(posedge clk)
begin
	if ((srst==1))
	hw <= 0;
  else if (clk_cycle_counter == 127)
  hw <= hw_read_in;
end

// rd_en_pulse: upon the 127th clock cycle of an episode we need a pulse to assert the start time of the (read from FIFOs and) send-out. here it is
always @ (posedge clk)
begin
if (srst==1)
rd_en_pulse <= 0;
else if (clk_cycle_counter==126)
rd_en_pulse <= 1;
else
rd_en_pulse <= 0;
end

// PC_out_temp: we need this signal to be decrement the weight of a read byte (in send-out phase) to zero in another register.
always @ (posedge clk)
begin
if (srst==1)	
PC_out_temp <= 0;	
else if (rd_en_pulse == 1)
PC_out_temp <= PC_out_temp; // just wait a cycle at the begining
else if ((PC_out_temp==0)&&(PC_out!=0))
PC_out_temp <= PC_out - 1;
else if (PC_out_temp==0)
PC_out_temp <= 0;
else
PC_out_temp <= PC_out_temp - 1;
end	

// The timing diagram below indicates why we need to infer PC_out_temp from PC_out in order to generate rd_en signals
// in fact, as previously stated, for 11001011 that has a weight of 5, five clock cycles are assigned, during which 
// rd_en is set only at the first cycle.

//##################EXAMPLE##################\\	
//#FIFO filled w/4 numbers whose weights are#\\
//#3,1,2, & 4. start signal is then asserted#\\
//###########################################\\
//#PC_out_temp#|0|0|0|0|2|1|0|0|1|0|3|2|1|0|#\\
//#PC_out######|X|X|X|3|3|3|1|2|2|4|4|4|4|0|#\\
//#rd_en#######|0|0|1|0|0|1|1|0|1|0|0|0|1|0|#\\
//#start_reg###|0|1|0|0|0|0|0|0|0|0|0|0|0|0|#\\
//#srst########|1|0|0|0|0|0|0|0|0|0|0|0|0|0|#\\
//###########################################\\


//Place holders: mutually exclusive pulses that are place holders for the outputs of the weight_locator. 
//A timing diagram of these signals are depicted at Wires and Registers section
always @ (posedge clk)
if (srst==1)
begin
L0_h<=0;
L1_h<=0;
L2_h<=0;
L3_h<=0;
L4_h<=0;
L5_h<=0;
L6_h<=0;
L7_h<=0;
end
else if (rd_en==1)
begin
L0_h<=1;
L1_h<=0;
L2_h<=0;
L3_h<=0;
L4_h<=0;
L5_h<=0;
L6_h<=0;
L7_h<=0;
end
else 
begin
L0_h<=0;
L1_h<=L0_h;
L2_h<=L1_h;
L3_h<=L2_h;
L4_h<=L3_h;
L5_h<=L4_h;
L6_h<=L5_h;
L7_h<=L6_h;
end


//this FIFO saves the non-zero bytes from input
fifo648 U1
       (
        .clk(clk) ,//input
        .srst(srst) ,//input
        .din(din_reg) ,//input
        .rd_en(rd_en) ,//input
        .wr_en(wr_en) ,//input
        .dout (stored_non_zero_byte) ,//output
        .full(overflow) ,//output, for future use
        .empty() //output, for future use
      );	   

//this FIFO saves the time (number of clock cycle in an episode) at which the non-zero byte was saved      
fifo648 U2
       (
        .clk(clk) ,//input
        .srst(srst) ,//input
        .din(clk_cycle_counter) ,//input
        .rd_en(rd_en) ,//input
        .wr_en(wr_en) ,//input
        .dout (stored_clk_cycle) ,//output
        .full() ,//output, for future use
        .empty() //output, for future use
      );	   

//This is the decoded, which is purely combinational. It generates the location of 1s in a byte on to its 8 index-outputs.
//meanwhile in generates the instant hamming weight of the given byte  
weight_locator U3 
		(
		.R(stored_non_zero_byte), //input
		.PC(PC_out), //output
		.L0(L0),//output
		.L1(L1),//output
		.L2(L2),//output
		.L3(L3),//output
		.L4(L4),//output
		.L5(L5),//output
		.L6(L6),//output
		.L7(L7)//output
		);

//    An Example to illustrate how the weight_locator works
//
//    |''''''''''''''''''|
//    |                PC|--5
// 1--|                L0|--0
// 1--|                L1|--1
// 0--|                L2|--4
// 0--|                L3|--6
// 1--|                L4|--7
// 0--|                L5|--0
// 1--|                L6|--0
// 1--|                L7|--0  
//    |..................|--0
//
// Note that in the above circuit PC=5 distinguishes 
// L0=0 as a 1-indicator from L5=0 as a non-1-indicator	 


// combining all  8 signals from weight_locator and 8 mutually exclusive pulses to represent the location of 1s at consecutive cycles
assign location_in_byte = L0_h*L0+L1_h*L1+L2_h*L2+L3_h*L3+L4_h*L4+L5_h*L5+L6_h*L6+L7_h*L7;
// calculating the location in 1028 bit stream based on the location at byte, and the clock cycle the byte came in
assign locations = location_in_byte+8*stored_clk_cycle;
// the span at which the outputs are valid 
assign valid = (valid_interval!=0);
// accumulating hamming weigh in read in phase
assign hw_read_in = PC_in + hw_reg;
// at send out phase we need to read from the FIFO at specific times, and not continuously.
assign rd_en_valid = (valid_interval!=0)&&(valid_interval!=1);
assign rd_en = (rd_en_pulse)||(((PC_out_temp==1)||(PC_out==1))&& rd_en_valid);
// at read in phase, if the input data is non-zero, signal wr_en will be set in order to have it stored
assign wr_en = (~start_reg) && (din_reg!=0) && (clk_cycle_counter<128);

endmodule